class dff_sequencer extends uvm_sequencer#(dff_seq_item);
  `uvm_component_utils(dff_sequencer) // reg class to uvm factory
  
  //standard constructor
  function new(string name ="dff_sequencer", uvm_component parent);
    super.new(name, parent);
    `uvm_info("sequencer Class", "constructor", UVM_MEDIUM)
  endfunction
  
  
endclass
